///////////////////////////////////////////////////
// HA.sv  This design will take in 3 bits       //
// and add them to produce a sum and carry out //
////////////////////////////////////////////////
module HA(
  input 	A,Cin,	// three input bits to be added
  output	S,Cout	 // Sum and carry out
);

	/////////////////////////////////////////////////
	// Declare any internal signals as type logic //
	///////////////////////////////////////////////

	/////////////////////////////////////////////////
	// Implement Full Adder as structural verilog //
	///////////////////////////////////////////////
	xor iXOR1(S,A,Cin);
	and iAND1(Cout,A,Cin);

endmodule
